library verilog;
use verilog.vl_types.all;
entity SHIFT_OPERATOR_vlg_sample_tst is
    port(
        \in\            : in     vl_logic_vector(3 downto 0);
        sleft           : in     vl_logic;
        sright          : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end SHIFT_OPERATOR_vlg_sample_tst;
