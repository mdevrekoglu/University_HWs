library verilog;
use verilog.vl_types.all;
entity ALU_2020510014_2020510028_2021510022_vlg_check_tst is
    port(
        overflow        : in     vl_logic;
        Rout            : in     vl_logic_vector(3 downto 0);
        sampler_rx      : in     vl_logic
    );
end ALU_2020510014_2020510028_2021510022_vlg_check_tst;
