library verilog;
use verilog.vl_types.all;
entity SHIFT_OPERATOR_vlg_vec_tst is
end SHIFT_OPERATOR_vlg_vec_tst;
